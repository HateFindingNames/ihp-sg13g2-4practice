** sch_path: /foss/designs/practicing/TempSensor/design_data/xschem/ptat_bjt_nmos-curr-mirror.sch
**.subckt ptat_bjt_nmos-curr-mirror
XM1 net1 net1 vh GND sg13_lv_nmos w=5u l=2u ng=1 m=1
XM2 VDD net1 vl GND sg13_lv_nmos w=5u l=2u ng=1 m=10
I1 GND net1 10u
Vgs2 VDD GND 1.2
XQ1 vh vh GND GND npn13G2 Nx=1
XQ2 vl vl GND GND npn13G2 Nx=1
**** begin user architecture code


.param temp 27
.control

save all
dc temp 0 100 1

let vdiff = vh - vl

wrdata ptat_bjt_nmos-curr-mirror.csv vdiff vh vl
write ptat_bjt_nmos-curr-mirror.raw

.endc




** IHP models
.lib cornerMOSlv.lib mos_tt
.lib cornerHBT.lib hbt_typ


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
