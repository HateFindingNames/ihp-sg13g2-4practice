** sch_path: /foss/designs/practicing/TempSensor/design_data/xschem/diff_amp_8-16_tb.sch
**.subckt diff_amp_8-16_tb
V2 inn GND 1m
V1 inp GND 10m
V3 net1 GND 1.263
x1 net1 inn inp out net2 diff_amp_8-16
XR1 GND out rhigh w=0.5e-6 l=5e-6 m=1 b=0
V4 net2 GND -1.263
**** begin user architecture code


** IHP models
.lib cornerMOSlv.lib mos_tt
.lib cornerCAP.lib cap_typ
.lib cornerRES.lib res_typ




.control

set tbname=diff_amp_8-16_tb
save dbgain gain out inp inn

dc V1 2m 200m 0.1m

let indiff = inp - inn
*if $out < 0
* let $out == 1e-12
*end
let gain = out / indiff
let dbgain = db(gain)

wrdata {$tbname}.csv gain out inp inn
write {$tbname}.raw

.endc


**** end user architecture code
**.ends

* expanding   symbol:  practicing/TempSensor/design_data/xschem/diff_amp_8-16.sym # of pins=5
** sym_path: /foss/designs/practicing/TempSensor/design_data/xschem/diff_amp_8-16.sym
** sch_path: /foss/designs/practicing/TempSensor/design_data/xschem/diff_amp_8-16.sch
.subckt diff_amp_8-16 vp inn inp out vn
*.ipin inp
*.opin out
*.ipin inn
*.iopin vn
*.iopin vp
XM6 net10 inn net2 vn sg13_lv_nmos w=10u l=0.5u ng=1 m=1
XM5 net11 inp net2 vn sg13_lv_nmos w=10u l=0.5u ng=1 m=1
XM2 net1 net1 net4 vp sg13_lv_pmos w=10u l=2u ng=1 m=10
XM1 net4 net1 vp vp sg13_lv_pmos w=6u l=1u ng=1 m=1
XM3 net3 net1 vp vp sg13_lv_pmos w=6u l=1u ng=1 m=1
XM4 net5 net1 net3 vp sg13_lv_pmos w=10u l=2u ng=1 m=10
XM7 net5 net5 net6 vn sg13_lv_nmos w=10u l=2u ng=1 m=10
XM8 net6 net5 vn vn sg13_lv_nmos w=10u l=5u ng=1 m=1
XM9 net2 net5 net7 vn sg13_lv_nmos w=10u l=2u ng=1 m=10
XM10 net7 net5 vn vn sg13_lv_nmos w=10u l=5u ng=1 m=1
XM15 net8 net8 vn vn sg13_lv_nmos w=10u l=1.5u ng=1 m=1
XM16 net9 net8 vn vn sg13_lv_nmos w=10u l=1.5u ng=1 m=1
XM11 net10 net1 vp vp sg13_lv_pmos w=10u l=1.67u ng=1 m=1
XM12 net8 net1 net10 vp sg13_lv_pmos w=10u l=2u ng=1 m=10
XM13 net11 net1 vp vp sg13_lv_pmos w=10u l=1.67u ng=1 m=1
XM14 net9 net1 net11 vp sg13_lv_pmos w=10u l=2u ng=1 m=10
XM17 out net1 vp vp sg13_lv_pmos w=9u l=5u ng=1 m=10
XM18 out net9 vn vn sg13_lv_nmos w=10u l=0.5u ng=1 m=5
I0 net1 vn 20u
XC2 out net9 cap_cmim w=35e-6 l=35e-6 m=1
.ends

.GLOBAL GND
.end
