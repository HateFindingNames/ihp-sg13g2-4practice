** sch_path: /foss/designs/practicing/TempSensor/design_data/xschem/device_testbenches/dc_res_temp.sch
**.subckt dc_res_temp
Vres Vcc GND 1.5
Vsil Vcc net1 0
.save i(vsil)
Vppd Vcc net2 0
.save i(vppd)
Vrh Vcc net3 0
.save i(vrh)
XR1 GND net1 rsil w=0.5e-6 l=1.5e-6 m=1 b=0
XR2 GND net2 rppd w=0.5e-6 l=0.5e-6 m=1 b=0
XR3 GND net3 rhigh w=0.5e-6 l=0.5e-6 m=1 b=0
**** begin user architecture code

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ_stat



.param temp=27
.control
save all
op
echo Silicide resisotr value:
print Vcc/I(Vsil)
echo Unsilicide poly resisotr value:
print Vcc/I(Vppd)
echo High poly resisotr value:
print Vcc/I(Vrh)
*reset
dc temp -40 125 1

let rrsil_perc = v(vcc)/(i(vsil)*38.59)
let rrppd_perc = v(vcc)/(i(vppd)*396.9)
let rrrh_perc = v(vcc)/(i(vrh)*1798)

let rrsil_abs = v(vcc)/i(vsil)
let rrppd_abs = v(vcc)/i(vppd)
let rrrh_abs = v(vcc)/i(vrh)

write dc_res_temp.raw
wrdata dc_res_temp.csv I(Vsil) I(Vppd) I(Vrh)
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
