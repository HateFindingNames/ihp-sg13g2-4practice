** sch_path: /foss/designs/practicing/TempSensor/design_data/xschem/ptat_nmos_only.sch
**.subckt ptat_nmos_only
XM1 Vdd net1 net1 GND sg13_lv_nmos w={inp_w} l={inp_l} ng=1 m=1
XM2 net1 net2 net2 GND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM3 net2 net3 net3 GND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM4 net3 GND GND GND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM5 Vdd net1 vout GND sg13_lv_nmos w={inp_w} l={inp_l} ng=1 m=1
XM7 Vdd net1 net4 GND sg13_lv_nmos w={inp_w} l={inp_l} ng=1 m=1
V1 Vdd GND 1
XM9 net5 net4 vout Vdd sg13_lv_pmos w={out_w} l={out_l} ng=1 m=1
XM6 GND net5 vout Vdd sg13_lv_pmos w={out_w} l={out_l} ng=1 m=1
**** begin user architecture code

.lib cornerMOSlv.lib mos_tt



.param inp_w = 0.15u inp_l = 0.13u
.param out_w = 0.15u out_l = 0.13u

.control

let run = 0
set curplot = new            ; 'new' creates a new plot of some name
set scratch = $curplot       ; the new plot is stored in 'scratch'
setplot $scratch

* Initialize a vector to store the results of each parameter alteration
let varinpl = unitvec(2)     ; Adjust the length according to the number of iterations

foreach varval 0.15u 0.3u
 alterparam inp_l = $varval
 echo '=== varval = $varval'
 dc temp 0 125 1
 set run = $&run
 let dt = $curplot            ; store the current plot name
 setplot $scratch             ; select the scratch plot
 let varinpl[$run] = $dt.vout ; Track results, indexed by the value being varied
 setplot $dt
 let run = run + 1
 reset
end

wrdata ptat_nmos_only_varinpl.csv {$scratch}.varinpl
write ptat_nmos_only_varinpl.raw

.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
