** sch_path: /foss/designs/practicing/TempSensor/design_data/xschem/a-210nW-npn-based-temp-sens.sch
**.subckt a-210nW-npn-based-temp-sens
XM1 net2 net2 vcc vcc sg13_lv_pmos w=5u l=2u ng=1 m=1
XM2 net3 net2 vcc vcc sg13_lv_pmos w=5u l=2u ng=1 m=10
XM3 vl net2 vcc vcc sg13_lv_pmos w=5u l=2u ng=1 m=1
XM4 vh net2 vcc vcc sg13_lv_pmos w=5u l=2u ng=1 m=1
XQ1 net2 net3 net1 net4 npn13G2 Nx=1
XQ2 net3 net3 GND net5 npn13G2 Nx=1
XQ3 vl vl GND net6 npn13G2 Nx=1
XQ4 vh vh GND net7 npn13G2 Nx=1
XR1 GND net1 rppd w=0.5e-6 l=0.5e-6 m=1 b=0
V1 vcc GND 1.5
**** begin user architecture code


.param temp 27
.control

save all
dc temp 0 100 1

let vdiff = vh - vl

wrdata ptat_bjt_nmos-curr-mirror.csv vdiff vh vl
write ptat_bjt_nmos-curr-mirror.raw

.endc




** IHP models
.lib cornerMOSlv.lib mos_tt
.lib cornerHBT.lib hbt_typ
.include ptat_bjt_nmos-curr-mirror.save


**** end user architecture code
**.ends
.GLOBAL GND
.end
