** sch_path: /foss/designs/practicing/TempSensor/design_data/xschem/diff_amp.sch
**.subckt diff_amp vdd v+ v- gnd out
*.ipin inp
*.opin out
*.ipin inn
*.iopin vn
*.iopin vp
*.ipin inp
*.ipin inn
XM6 net10 inn net2 vn sg13_lv_nmos w=10u l=0.5u ng=1 m=1
XM5 net11 inp net2 vn sg13_lv_nmos w=10u l=0.5u ng=1 m=1
XM2 net12 net1 net4 vp sg13_lv_pmos w=10u l=2u ng=1 m=10
XM1 net4 net1 vp vp sg13_lv_pmos w=6u l=1u ng=1 m=1
XM3 net3 net1 vp vp sg13_lv_pmos w=6u l=1u ng=1 m=1
XM4 net5 net1 net3 vp sg13_lv_pmos w=10u l=2u ng=1 m=10
XM7 net5 net5 net6 vn sg13_lv_nmos w=10u l=2u ng=1 m=10
XM8 net6 net5 vn vn sg13_lv_nmos w=10u l=5u ng=1 m=1
XM9 net2 net5 net7 vn sg13_lv_nmos w=10u l=2u ng=1 m=10
XM10 net7 net5 vn vn sg13_lv_nmos w=10u l=5u ng=1 m=1
XM15 net8 net8 vn vn sg13_lv_nmos w=10u l=1.5u ng=1 m=1
XM16 net9 net8 vn vn sg13_lv_nmos w=10u l=1.5u ng=1 m=1
XM11 net10 net1 vp vp sg13_lv_pmos w=10u l=1.67u ng=1 m=1
XM12 net8 net1 net10 vp sg13_lv_pmos w=10u l=2u ng=1 m=10
XM13 net11 net1 vp vp sg13_lv_pmos w=10u l=1.67u ng=1 m=1
XM14 net9 net1 net11 vp sg13_lv_pmos w=10u l=2u ng=1 m=10
XM17 out net1 vp net13 sg13_lv_pmos w=9u l=5u ng=1 m=10
XM18 out net9 vn vn sg13_lv_nmos w=10u l=0.5u ng=1 m=5
I0 net12 vn 20u
XC2 net9 out cap_cmim w=35e-6 l=35e-6 m=1
V1 inp GND 10.1m
V2 inn GND 10m
**** begin user architecture code


** IHP models
.lib cornerMOSlv.lib mos_tt
.lib cornerCAP.lib cap_typ




.param temp 27
.control

set tbname=op-amp_1
save all
dc in+ 10m 12m 0.01m

let vdiff = inp - inn

wrdata {$tbname}.csv vdiff out inp inn
write {$tbname}.raw

.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
