** sch_path: /foss/designs/practicing/TempSensor/design_data/xschem/snoa748c_temp_sensor_tb.sch
**.subckt snoa748c_temp_sensor_tb
XQ1 net1 net1 GND GND npn13G2 Nx=1
XQ2 vl net1 net2 net2 npn13G2 Nx=1
I0 GND net1 50u
V1 vh GND 1.2
XR1 GND net2 rppd w=0.5e-6 l=0.5e-6 m=1 b=0
XR2 vl vh rppd w=0.5e-6 l=0.5e-6 m=1 b=0
**** begin user architecture code


.param temp 27
.control

save all
dc temp 0 100 1

let vdiff = vl - vh

wrdata ptat_bjt_nmos-curr-mirror.csv vdiff vh vl
write ptat_bjt_nmos-curr-mirror.raw

.endc




** IHP models
.lib cornerRES.lib res_typ
.lib cornerHBT.lib hbt_typ


**** end user architecture code
**.ends
.GLOBAL GND
.end
