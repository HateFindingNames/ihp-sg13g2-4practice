** sch_path: /foss/designs/practicing/TempSensor/design_data/xschem/diff_amp_test.sch
**.subckt diff_amp_test
XM2 net2 net1 net1 net2 sg13_lv_nmos w=7.0u l=1u ng=1 m=1
XM1 out net5 net3 GND sg13_lv_nmos w=0.35u l=10u ng=1 m=1
XM3 net2 net1 out net2 sg13_lv_nmos w=7.0u l=1u ng=1 m=1
XM4 net1 net4 net3 GND sg13_lv_nmos w=1.0u l=10u ng=1 m=1
XM5 net3 net2 GND GND sg13_lv_nmos w=1.0u l=1u ng=1 m=1
V1 net4 GND 100m
V2 net5 GND 2
V3 net2 GND 2
**** begin user architecture code


.temp 27
.control
save all
dc V2 100m 150m 10u
write diff_amp_test.raw
.endc




** IHP models
.lib cornerMOSlv.lib mos_tt


**** end user architecture code
**.ends
.GLOBAL GND
.end
